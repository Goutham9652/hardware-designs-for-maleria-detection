
`timescale 1ns / 1ps

module cnn_top_tb;
    // Parameters (using smaller values for simulation)
    parameter INPUT_SIZE = 64;  // Using 16x16 for testing
    parameter KERNEL_SIZE = 3;
    parameter CONV_OUTPUT_SIZE = INPUT_SIZE - KERNEL_SIZE + 1;    // 14
    parameter PAD_OUTPUT_SIZE = CONV_OUTPUT_SIZE + 2;            // 16
    parameter POOL_OUTPUT_SIZE = PAD_OUTPUT_SIZE / 2;            // 8
    
    // Bit width calculations
    parameter INPUT_BITS = INPUT_SIZE * INPUT_SIZE;
    parameter CONV_OUTPUT_BITS = CONV_OUTPUT_SIZE * CONV_OUTPUT_SIZE * 4;
    parameter PAD_OUTPUT_BITS = PAD_OUTPUT_SIZE * PAD_OUTPUT_SIZE * 4;
    parameter POOL_OUTPUT_BITS = POOL_OUTPUT_SIZE * POOL_OUTPUT_SIZE * 4;
    
    // Test bench signals
    reg clk;
    reg rst;
    reg start;
    reg [INPUT_BITS-1:0] input_image;
    wire result;
    wire done;
    
    // Internal probes for debugging
    wire [CONV_OUTPUT_BITS-1:0] conv_output;
    wire [PAD_OUTPUT_BITS-1:0] pad_output;
    wire [POOL_OUTPUT_BITS-1:0] pool_output;
    wire conv_done, pad_done, pool_done, classify_done;
    
    // DUT Instantiation
    cnn_top #(
        .INPUT_SIZE(INPUT_SIZE),
        .KERNEL_SIZE(KERNEL_SIZE)
    ) dut (
        .clk(clk),
        .rst(rst),
        .start(start),
        .input_image(input_image),
        .result(result),
        .done(done)
    );
    
    // Connect internal signals for monitoring
    assign conv_output = dut.conv_output;
    assign pad_output = dut.pad_output;
    assign pool_output = dut.pool_output;
    assign conv_done = dut.conv_done;
    assign pad_done = dut.pad_done;
    assign pool_done = dut.pool_done;
    assign classify_done = dut.classify_done;
    
    // Clock generation
    initial begin
        clk = 0;
        forever #5 clk = ~clk;  // 100MHz clock
    end
    
    // Display the input image
    task display_input_image;
        integer i, j, idx;
        begin
            $display("\n===== INPUT IMAGE (%0d x %0d) =====", INPUT_SIZE, INPUT_SIZE);
            for (i = 0; i < INPUT_SIZE; i = i + 1) begin
                for (j = 0; j < INPUT_SIZE; j = j + 1) begin
                    idx = i * INPUT_SIZE + j;
                    $write("%b", input_image[idx]);
                end
                $write("\n");
            end
        end
    endtask
    
    // Display convolution output
    task display_conv_output;
        integer i, j, idx;
        reg [3:0] pixel;
        begin
            $display("\n===== CONVOLUTION OUTPUT (%0d x %0d) =====", CONV_OUTPUT_SIZE, CONV_OUTPUT_SIZE);
            for (i = 0; i < CONV_OUTPUT_SIZE; i = i + 1) begin
                for (j = 0; j < CONV_OUTPUT_SIZE; j = j + 1) begin
                    idx = (i * CONV_OUTPUT_SIZE + j) * 4;
                    pixel = conv_output[idx+:4]; // Extract 4 bits
                    $write("%d", pixel);
                end
                $write("\n");
            end
        end
    endtask
    
    // Display padding output
    task display_pad_output;
        integer i, j, idx;
        reg [3:0] pixel;
        begin
            $display("\n===== PADDING OUTPUT (%0d x %0d) =====", PAD_OUTPUT_SIZE, PAD_OUTPUT_SIZE);
            for (i = 0; i < PAD_OUTPUT_SIZE; i = i + 1) begin
                for (j = 0; j < PAD_OUTPUT_SIZE; j = j + 1) begin
                    idx = (i * PAD_OUTPUT_SIZE + j) * 4;
                    pixel = pad_output[idx+:4]; // Extract 4 bits
                    $write("%d", pixel);
                end
                $write("\n");
            end
        end
    endtask
    
    // Display pooling output
    task display_pool_output;
        integer i, j, idx;
        reg [3:0] pixel;
        begin
            $display("\n===== POOLING OUTPUT (%0d x %0d) =====", POOL_OUTPUT_SIZE, POOL_OUTPUT_SIZE);
            for (i = 0; i < POOL_OUTPUT_SIZE; i = i + 1) begin
                for (j = 0; j < POOL_OUTPUT_SIZE; j = j + 1) begin
                    idx = (i * POOL_OUTPUT_SIZE + j) * 4;
                    pixel = pool_output[idx+:4]; // Extract 4 bits
                    $write("%d", pixel);
                end
                $write("\n");
            end
        end
    endtask
    
    // Test stimulus
    initial begin
        // Initialize signals
        rst = 1;
        start = 0;
        input_image = 0;
        
        // Apply reset
        #20;
        rst = 0;
        #20;
        
        // Load test image (16x16 binary image)
        // Checkerboard pattern for testing
//        input_image = 256'b0000011000000000000111111100000000111111111100000111111111111000011111111111110011111111111111101111111111111111011111111111111101111111111111110111111111111111001111111111111100111111111111110001111111111110000001111111111000000111111111000000000011110000;
       // input_image = 64'b0000010001111110010011100100101100110010110001100111100000110000;
       //  input_image = 1024'b0000000000000011111000000000000000000000000011111111100000000000000000000111111111111111000000000000000011111111111111111000000000000011111111111111111111100000000000111111111111111111111000000000111111111111111111111111000000001111111111111111111111111000001111111111111111111111111110000011111111111111111111111111100001111111111111111111111111111100111111111111111111111111100111101111111111111111111111111001111001111111111111111111111111111111111111111111110011111110111111110111111111111110011111101111111101111111001111111111111111111111011111110001111111111111111111110111111100011111011111111111111100111111000011000011111111111111001111111000100000111111111111100011111111111000001111111111111000011111111111000111111111111110000110111111111111111111111111100001111111111111111111111111110000011111111111111111111111111000000011111111111111110111111110000000001111111111111101111111000000000001111111111111111111100000000000001111111111111111110000000000000000001111111111111000000000000000000000001111011000000000;
        input_image = 4096'b0000000000000000000000000111000000000000000000000000000000000000000000000000000000000000111111111110000000000000000000000000000000000000000000000000000111111111111000000000000000000000000000000000000000000000011111111111111111111110011110000000000000000000000000000000001111111111111111111111111111111100000000000000000000000000000000111111111111111111111111111111111000000000000000000000000000000111111111111111111111111111111111110000000000000000000000000000111111111111111111111111111111111111100000000000000000000000001111111111111111111111111111111111111111000000000000000000000011111111111111111111111111111111111111111110000000000000000000011111111111111111111111111111111111111111111110000000000000000011111111111111111111111111111111111111111111111000000000000000011111111111111111111111111111111111111111111111100000000000000011111111111111111111111111111111111111111111111111000000000000001111111111111111111111111111111111111111111111111110000000000000111111111111111111111111111111111111111111111111111110000000000011111111111111111111111111111111111111111111111111111000000000011111111111111111111111111111111111111111111111111111110000000001111111111111111111111111111111111111111111111111111111110000000111111111111111111111111111111111111111111111111111111111000000111111111111111111111111111111111111111111111111111111111110000011111111111111111111111111111111111111111111111111111111111000001111111111111111111111111111111111111111111111111111111111110011111111111111111111111111111111111111111111111111111111111111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001111111111111111111111111111111111111111111111111111111111111100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001111111111111111111111111111111111111111111111111111111111111000011111111111111111111111111111111111111111111111111111111111100001111111111111111111111111111111111111111111111111111111111110000011111111111111111111111111111111111111111111111111111111111000001111111111111111111111111111111111111111111111111111111111000000111111111111111111111111111111111111111111111111111111111100000011111111111111111111111111111111111111111111111111111111110000000111111111111111111111111111111111111111111111111111111111000000000111111111111111111111111111111111111111111111111111111100000000011111111111111111111111111111111111111111111111111111100000000001111111111111111111111111111111111111111111111111111100000000000011111111111111111111111111111111111111111111111111100000000000000111111111111111111111111111111111111111111111111100000000000000000111111111111111111111111111111111111111111111100000000000000000001111111111111111111111111111111111111111111100000000000000000000111111111111111111111111111111111111111111100000000000000000000000111111111111111111111111111111111111111100000000000000000000000001111111111111111111111111111111111111000000000000000000000000000011111111111111111111111111111111111000000000000000000000000000000111111111111111111111111111111111100000000000000000000000000000001111111111111111111111111111111100000000000000000000000000000000001111111111111111111111111110000000000000000000000000000000000000001111111111111111111111000000000000000000000000000000000000000000011111111111111111111000000000000000000000000000000000000000000000111111111111111111000000000000000000000000000000000000000000000000011100000000000000000000000000000000000;
        
        
        display_input_image();
        
        // Start processing
        #10;
        $display("Starting CNN processing at time %0t", $time);
        start = 1;
        
        // Wait for convolution to complete
        @(posedge conv_done);
        #10; // Wait for a few cycles for stability
        display_conv_output();
        
        // Wait for padding to complete
        @(posedge pad_done);
        #10; // Wait for a few cycles for stability
        display_pad_output();
        
        // Wait for pooling to complete
        @(posedge pool_done);
        #10; // Wait for a few cycles for stability
        display_pool_output();
        
        // Wait for done signal
        @(posedge done);
        $display("CNN processing completed at time %0t", $time);
        $display("Classification result: %s", result ? "Diseased" : "Healthy");
        
        // De-assert start and wait
        #20;
        start = 0;
        #50;
        
        // Allow simulation to complete
        #200;
        $display("Simulation completed at time %0t", $time);
        $finish;
    end
    
    // Monitor state transitions
    reg [2:0] prev_state;
    initial begin
        prev_state = 0;
        forever begin
            @(posedge clk);
            if (dut.state !== prev_state) begin
                case (dut.state)
                    0: $display("Time %0t: State -> IDLE", $time);
                    1: $display("Time %0t: State -> CONV_STAGE", $time);
                    2: $display("Time %0t: State -> PADDING_STAGE", $time);
                    3: $display("Time %0t: State -> POOLING_STAGE", $time);
                    4: $display("Time %0t: State -> CLASSIFY_STAGE", $time);
                    5: $display("Time %0t: State -> FINISHED", $time);
                    default: $display("Time %0t: State -> UNKNOWN (%0d)", $time, dut.state);
                endcase
                prev_state = dut.state;
            end
        end
    end
    
    // Monitor stage completion events
    initial begin
        forever begin
            @(posedge clk);
            if (conv_done && dut.state == 1)
                $display("Time %0t: Convolution stage completed", $time);
            if (pad_done && dut.state == 2)
                $display("Time %0t: Padding stage completed", $time);
            if (pool_done && dut.state == 3)
                $display("Time %0t: Pooling stage completed", $time);
            if (classify_done && dut.state == 4)
                $display("Time %0t: Classification stage completed", $time);
        end
    end
    
   
    
endmodule
